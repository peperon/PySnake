[DEFAULT]
level = 0
snake = [(48, 64), (64, 64)]
food = (546, 128)
direction = 4

